LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.EE232.ALL;

ENTITY DEMUX_1X2 IS

	PORT(X0, S: IN STD_LOGIC;
	Y0, Y1 : OUT STD_LOGIC);
END DEMUX_1X2;

ARCHITECTURE STRUCTURE OF DEMUX_1X2 IS
SIGNAL S0 : STD_LOGIC;

BEGIN
U0 : AND_2 port map (X0, S0, Y0);
U1 : NOT_1 port map(S, S0);
U2 : AND_2 port map (X0, S, Y1);


END STRUCTURE;
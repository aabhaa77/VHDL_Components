LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.EE232.ALL;

ENTITY DEMUX_1X4 IS

	PORT(I0: IN STD_LOGIC;
		S : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		O : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END DEMUX_1X4;


ARCHITECTURE STRUCTURE OF DEMUX_1X4 IS
SIGNAL Y0, Y1 : STD_LOGIC;

BEGIN
U0 : DEMUX_1X2 port map (I0, S(0), Y0, Y1);
U1 : DEMUX_1X2 port map(Y0, S(1), O(0), O(2));
U2 : DEMUX_1X2 port map(Y1, S(1), O(1), O(3));



END STRUCTURE;
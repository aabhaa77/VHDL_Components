LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.EE232.ALL;

ENTITY MUX_4X1 IS

	PORT(X0, X1, X2, X3, S0, S1: IN STD_LOGIC;
	Y : OUT STD_LOGIC);
END MUX_4X1;

ARCHITECTURE STRUCTURE OF MUX_4X1 IS
SIGNAL P0, P1 : STD_LOGIC;

BEGIN
U0 : MUX_2X1 port map (X0, S0, X1, P0);
U1 : MUX_2X1 port map(X2, S0, X3, P1);
U2 : MUX_2X1 port map (P0, S1, P1, Y);

END STRUCTURE;